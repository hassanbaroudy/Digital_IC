package pack1;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "hassan_sequence_item.sv"
`include "hassan_sequence.sv"
`include "hassan_driver.sv"
`include "hassan_monitor.sv"
`include "hassan_sequencer.sv"
`include "hassan_agent.sv"
`include "hassan_scoreboard.sv"
`include "hassan_subscriber.sv"
`include "hassan_env.sv"
`include "hassan_test.sv"
endpackage